library ieee;
use ieee.std_logic_1164.all;

entity jk_flip_flop is
    port (
        j, k, clk, reset: in std_logic;
        q, q_bar: out std_logic
    );
end entity jk_flip_flop;

architecture structural of jk_flip_flop is
    
end architecture structural;
